library verilog;
use verilog.vl_types.all;
entity problem_set2_schematic_vlg_vec_tst is
end problem_set2_schematic_vlg_vec_tst;
